package datatypes;
import FixedPoint::*;
 
typedef FixedPoint#(14,2) DataType;
typedef FixedPoint#(2,14) CoeffType;
typedef UInt#(16) BramWidth;
typedef UInt#(6) BramLength;

endpackage
