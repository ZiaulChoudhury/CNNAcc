package datatypes;
import FixedPoint::*;

`define IMG 8
#define Mr 1024

typedef FixedPoint#(10,6) DataType;
typedef FixedPoint#(2,14) CoeffType;
typedef UInt#(14) BramWidth;
typedef UInt#(6) BramLength;

endpackage
